header.welcome = välkommen
header.register = registrera
header.login = logga in
header.userview = applikant

title.index = cv registrering
title.register = registrera ny användare
title.login = logga in
title.userview = applikant
title.competence = lägg till ny kompetens
title.error = ett fel har inträffat 

error.competenceProfileNotFound = den valda kompetensprofilen hittades inte
error.competenceProfileNotYours = du kan inte ta bort kompetensprofiler du inte äger
error.availabilityNotFound = den valda tillgängligheten hittades inte
error.availabilityNotYours = du kan inte ta bort andra användares tillgänglighet
error.notAuthorized = endast rekryterare kan besöka denna sida
error.specComp = välj en kompetens

error.userNotFound = den valda användaren hittades inte
error.dateFormat = fel datumformat angivet
error.notfound = sidan hittades inte

userlist.users = Användare

button.login = logga in
button.logout = logga ut
button.register = registrera
button.registernew = registrera ny användare
button.addCompetence = lägg till kompetens
button.remove = ta bort
button.hire = anställ
button.deny = avslå
button.pdf = ladda ner pdf


change = ändra
save = spara

from = från
to = till

availability = tillgänglighet

panel.competenceName = typ av kompetens
panel.competenceYears = år av erfarenhet

plain.competence = kompetens

list.competences = kompetenser:

plain.username = användarnamn
choose.username = välj användarnamn

choose.password = välj lösenord
plain.password = lösenord
choose.confirmPassword = skriv in lösenordet igen
plain.confirmPassword = upprepa lösenord
choose.email = välj epostadress
plain.email = epostadress
choose.name = välj ditt förnamn
plain.name = förnamn
choose.surname = välj ditt efternamn
plain.surname = efternamn
choose.ssn = välj ditt personnummer
plain.ssn = personnummer
choose.competence = välj en kompetens

competence.1 = Projektledning
competence.2 = Multimediedesign
competence.3 = Korvgrillning
competence.4 = Karuselldrift


constraints.required = Obligatorisk

user.isHired = Du har blivit anställd!
user.notHiredYet = Du har inte blivit anställd än

password.length = lösenordet måste vara minst 6 tecken långt
