header.welcome = välkommen
header.register = registrera
header.login = logga in

title.index = cv registrering
title.register = registrera ny användare
title.login = logga in
title.competence = lägg till ny kompetens

button.login = logga in
button.logout = logga ut
button.register = registrera
button.registernew = registrera ny användare
button.addCompetence = lägg till kompetens

panel.competenceName = typ av kompetens
panel.competenceYears = år av erfarenhet

plain.competence = kompetens

list.competences = kompetenser:

choose.competence = välj en kompetens

competence.1 = korvgrillning
competence.2 = karusellåkning


