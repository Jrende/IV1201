header.welcome = välkommen
header.register = registrera
header.login = logga in

title.index = cv registrering
title.register = registrera ny användare
title.login = logga in

button.login = logga in
button.logout = logga ut
button.register = registrera
button.registernew = registrera ny användare